`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:50:38 10/17/2022 
// Design Name: 
// Module Name:    lab5_1017_verilog 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab5_1017_verilog(
    input A,
    input B,
    input C,
    input D,
    input S0,
    input S1,
    input S2,
    output Y
    );


endmodule
